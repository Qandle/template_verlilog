module light (
    output led
);
    assign led = 1'b1;
endmodule
